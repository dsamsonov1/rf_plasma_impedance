.title KiCad schematic
R2 5 4 0.5
V0 1 0 SINE(0 100 13.56e6 0 0)
R1 2 1 50
L1 4 3 1.237u
C1 2 0 1.249n
R3 6 0 0.5
C5 2 3 166p
B1 5 7 i=v(7,5) > 0 ? 2.914584967225386*exp(-0.2105951039219109*v(7,5)) : 1e-12
I2 9 10 0.020305703373389043
C4 9 10 C='sqrt(7.965e-19/abs(v(9,10)))'
L2 8 7 162.272n
R4 9 8 9.72264147439682
B2 10 9 i=v(9,10) > 0 ? 8.743754901676157*exp(-0.2105951039219109*v(9,10)) : 1e-12
V1 10 0 0
I1 7 5 0.006768567791129681
C2 6 5 200p
C3 7 5 C='sqrt(8.85e-20/abs(v(7,5)))'
.end
